-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Sat Feb 08 19:57:21 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY mdr IS 
	PORT
	(	
		clk :  IN  STD_LOGIC;
		clear :  IN  STD_LOGIC;
		MDRin :  IN  STD_LOGIC;
		Read :  IN  STD_LOGIC;
		BusMuxOut :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		MemDataIn :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		MDRDataOut :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END mdr;

ARCHITECTURE bdf_type OF mdr IS 

COMPONENT mux2to1_32
	PORT(SEL : IN STD_LOGIC;
		 X0_in : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 X1_in : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Y : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT reg32
	PORT(clk : IN STD_LOGIC;
		 reset_n : IN STD_LOGIC;
		 en : IN STD_LOGIC;
		 d : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN

b2v_read_select : mux2to1_32
PORT MAP(SEL => Read,
		 X0_in => BusMuxOut,
		 X1_in => MemDataIn,
		 Y => SYNTHESIZED_WIRE_0);

b2v_mdr_reg : reg32
PORT MAP(clk => clk,
		 reset_n => clear,
		 en => MDRin,
		 d => SYNTHESIZED_WIRE_0,
		 q => MDRDataOut);


END bdf_type;